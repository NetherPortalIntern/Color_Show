library verilog;
use verilog.vl_types.all;
entity tb_config is
end tb_config;
