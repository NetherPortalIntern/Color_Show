library verilog;
use verilog.vl_types.all;
entity tb_Counter is
end tb_Counter;
