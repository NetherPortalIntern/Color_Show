library verilog;
use verilog.vl_types.all;
entity tb_Clock_Divider is
end tb_Clock_Divider;
