library verilog;
use verilog.vl_types.all;
entity tb_DB is
end tb_DB;
